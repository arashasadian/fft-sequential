library ieee;
use ieee.std_logic_1164.all;

package fftpackage is

    type array_of_integer is array(natural range <>) of integer;
    type array_2d is array(natural range <>) of array_of_integer;

    constant SIZE : integer := 8;
    constant rom_shift_amount : integer := -4;
    signal sin_rom, cos_rom : array_of_integer(360 downto 0);
    procedure rom_generator(signal enable : in std_logic; signal s_rom, c_rom : inout array_of_integer(360 downto 0));

    component fft2 is
        generic (rows, cols : integer := SIZE);
        port(
            input_array : in array_2d(rows - 1 downto 0)(cols - 1 downto 0);
            output_array_real : out array_2d(rows - 1 downto 0)(cols - 1 downto 0);
            output_array_imag : out array_2d(rows - 1 downto 0)(cols - 1 downto 0)
        );
    end component fft2;

    component fft is
        generic (size : integer := SIZE);
        port (clk :in std_logic;
            input_array : in array_of_integer(size - 1 downto 0);
            input_array_imag : in array_of_integer(size-1 downto 0);
            output_real_array, output_imag_array : out array_of_integer(size - 1 downto 0);
            end_sig : out std_logic
        );
    end component fft;

    component dft is
        generic (size : integer := SIZE/2);
        port (clk :in std_logic;
            input_array_real : in array_of_integer(size - 1 downto 0);
            input_array_imag : in array_of_integer(size - 1 downto 0);
            output_real_array, output_imag_array : out array_of_integer(size - 1 downto 0);
            done : out std_logic
        );
    end component dft;
    

end package fftpackage;

package body fftpackage is

    procedure rom_generator (signal enable : in std_logic; 
        signal s_rom, c_rom : inout array_of_integer(360 downto 0)) is
        begin
            if rising_edge(enable) then
                s_rom(0) <= 0;
s_rom(1) <= 17;
s_rom(2) <= 34;
s_rom(3) <= 52;
s_rom(4) <= 69;
s_rom(5) <= 87;
s_rom(6) <= 104;
s_rom(7) <= 121;
s_rom(8) <= 139;
s_rom(9) <= 156;
s_rom(10) <= 173;
s_rom(11) <= 190;
s_rom(12) <= 207;
s_rom(13) <= 224;
s_rom(14) <= 241;
s_rom(15) <= 258;
s_rom(16) <= 275;
s_rom(17) <= 292;
s_rom(18) <= 309;
s_rom(19) <= 325;
s_rom(20) <= 342;
s_rom(21) <= 358;
s_rom(22) <= 374;
s_rom(23) <= 390;
s_rom(24) <= 406;
s_rom(25) <= 422;
s_rom(26) <= 438;
s_rom(27) <= 453;
s_rom(28) <= 469;
s_rom(29) <= 484;
s_rom(30) <= 499;
s_rom(31) <= 515;
s_rom(32) <= 529;
s_rom(33) <= 544;
s_rom(34) <= 559;
s_rom(35) <= 573;
s_rom(36) <= 587;
s_rom(37) <= 601;
s_rom(38) <= 615;
s_rom(39) <= 629;
s_rom(40) <= 642;
s_rom(41) <= 656;
s_rom(42) <= 669;
s_rom(43) <= 681;
s_rom(44) <= 694;
s_rom(45) <= 707;
s_rom(46) <= 719;
s_rom(47) <= 731;
s_rom(48) <= 743;
s_rom(49) <= 754;
s_rom(50) <= 766;
s_rom(51) <= 777;
s_rom(52) <= 788;
s_rom(53) <= 798;
s_rom(54) <= 809;
s_rom(55) <= 819;
s_rom(56) <= 829;
s_rom(57) <= 838;
s_rom(58) <= 848;
s_rom(59) <= 857;
s_rom(60) <= 866;
s_rom(61) <= 874;
s_rom(62) <= 882;
s_rom(63) <= 891;
s_rom(64) <= 898;
s_rom(65) <= 906;
s_rom(66) <= 913;
s_rom(67) <= 920;
s_rom(68) <= 927;
s_rom(69) <= 933;
s_rom(70) <= 939;
s_rom(71) <= 945;
s_rom(72) <= 951;
s_rom(73) <= 956;
s_rom(74) <= 961;
s_rom(75) <= 965;
s_rom(76) <= 970;
s_rom(77) <= 974;
s_rom(78) <= 978;
s_rom(79) <= 981;
s_rom(80) <= 984;
s_rom(81) <= 987;
s_rom(82) <= 990;
s_rom(83) <= 992;
s_rom(84) <= 994;
s_rom(85) <= 996;
s_rom(86) <= 997;
s_rom(87) <= 998;
s_rom(88) <= 999;
s_rom(89) <= 999;
s_rom(90) <= 1000;
s_rom(91) <= 999;
s_rom(92) <= 999;
s_rom(93) <= 998;
s_rom(94) <= 997;
s_rom(95) <= 996;
s_rom(96) <= 994;
s_rom(97) <= 992;
s_rom(98) <= 990;
s_rom(99) <= 987;
s_rom(100) <= 984;
s_rom(101) <= 981;
s_rom(102) <= 978;
s_rom(103) <= 974;
s_rom(104) <= 970;
s_rom(105) <= 965;
s_rom(106) <= 961;
s_rom(107) <= 956;
s_rom(108) <= 951;
s_rom(109) <= 945;
s_rom(110) <= 939;
s_rom(111) <= 933;
s_rom(112) <= 927;
s_rom(113) <= 920;
s_rom(114) <= 913;
s_rom(115) <= 906;
s_rom(116) <= 898;
s_rom(117) <= 891;
s_rom(118) <= 882;
s_rom(119) <= 874;
s_rom(120) <= 866;
s_rom(121) <= 857;
s_rom(122) <= 848;
s_rom(123) <= 838;
s_rom(124) <= 829;
s_rom(125) <= 819;
s_rom(126) <= 809;
s_rom(127) <= 798;
s_rom(128) <= 788;
s_rom(129) <= 777;
s_rom(130) <= 766;
s_rom(131) <= 754;
s_rom(132) <= 743;
s_rom(133) <= 731;
s_rom(134) <= 719;
s_rom(135) <= 707;
s_rom(136) <= 694;
s_rom(137) <= 681;
s_rom(138) <= 669;
s_rom(139) <= 656;
s_rom(140) <= 642;
s_rom(141) <= 629;
s_rom(142) <= 615;
s_rom(143) <= 601;
s_rom(144) <= 587;
s_rom(145) <= 573;
s_rom(146) <= 559;
s_rom(147) <= 544;
s_rom(148) <= 529;
s_rom(149) <= 515;
s_rom(150) <= 499;
s_rom(151) <= 484;
s_rom(152) <= 469;
s_rom(153) <= 453;
s_rom(154) <= 438;
s_rom(155) <= 422;
s_rom(156) <= 406;
s_rom(157) <= 390;
s_rom(158) <= 374;
s_rom(159) <= 358;
s_rom(160) <= 342;
s_rom(161) <= 325;
s_rom(162) <= 309;
s_rom(163) <= 292;
s_rom(164) <= 275;
s_rom(165) <= 258;
s_rom(166) <= 241;
s_rom(167) <= 224;
s_rom(168) <= 207;
s_rom(169) <= 190;
s_rom(170) <= 173;
s_rom(171) <= 156;
s_rom(172) <= 139;
s_rom(173) <= 121;
s_rom(174) <= 104;
s_rom(175) <= 87;
s_rom(176) <= 69;
s_rom(177) <= 52;
s_rom(178) <= 34;
s_rom(179) <= 17;
s_rom(180) <= 0;
s_rom(181) <= -17;
s_rom(182) <= -34;
s_rom(183) <= -52;
s_rom(184) <= -69;
s_rom(185) <= -87;
s_rom(186) <= -104;
s_rom(187) <= -121;
s_rom(188) <= -139;
s_rom(189) <= -156;
s_rom(190) <= -173;
s_rom(191) <= -190;
s_rom(192) <= -207;
s_rom(193) <= -224;
s_rom(194) <= -241;
s_rom(195) <= -258;
s_rom(196) <= -275;
s_rom(197) <= -292;
s_rom(198) <= -309;
s_rom(199) <= -325;
s_rom(200) <= -342;
s_rom(201) <= -358;
s_rom(202) <= -374;
s_rom(203) <= -390;
s_rom(204) <= -406;
s_rom(205) <= -422;
s_rom(206) <= -438;
s_rom(207) <= -453;
s_rom(208) <= -469;
s_rom(209) <= -484;
s_rom(210) <= -500;
s_rom(211) <= -515;
s_rom(212) <= -529;
s_rom(213) <= -544;
s_rom(214) <= -559;
s_rom(215) <= -573;
s_rom(216) <= -587;
s_rom(217) <= -601;
s_rom(218) <= -615;
s_rom(219) <= -629;
s_rom(220) <= -642;
s_rom(221) <= -656;
s_rom(222) <= -669;
s_rom(223) <= -681;
s_rom(224) <= -694;
s_rom(225) <= -707;
s_rom(226) <= -719;
s_rom(227) <= -731;
s_rom(228) <= -743;
s_rom(229) <= -754;
s_rom(230) <= -766;
s_rom(231) <= -777;
s_rom(232) <= -788;
s_rom(233) <= -798;
s_rom(234) <= -809;
s_rom(235) <= -819;
s_rom(236) <= -829;
s_rom(237) <= -838;
s_rom(238) <= -848;
s_rom(239) <= -857;
s_rom(240) <= -866;
s_rom(241) <= -874;
s_rom(242) <= -882;
s_rom(243) <= -891;
s_rom(244) <= -898;
s_rom(245) <= -906;
s_rom(246) <= -913;
s_rom(247) <= -920;
s_rom(248) <= -927;
s_rom(249) <= -933;
s_rom(250) <= -939;
s_rom(251) <= -945;
s_rom(252) <= -951;
s_rom(253) <= -956;
s_rom(254) <= -961;
s_rom(255) <= -965;
s_rom(256) <= -970;
s_rom(257) <= -974;
s_rom(258) <= -978;
s_rom(259) <= -981;
s_rom(260) <= -984;
s_rom(261) <= -987;
s_rom(262) <= -990;
s_rom(263) <= -992;
s_rom(264) <= -994;
s_rom(265) <= -996;
s_rom(266) <= -997;
s_rom(267) <= -998;
s_rom(268) <= -999;
s_rom(269) <= -999;
s_rom(270) <= -1000;
s_rom(271) <= -999;
s_rom(272) <= -999;
s_rom(273) <= -998;
s_rom(274) <= -997;
s_rom(275) <= -996;
s_rom(276) <= -994;
s_rom(277) <= -992;
s_rom(278) <= -990;
s_rom(279) <= -987;
s_rom(280) <= -984;
s_rom(281) <= -981;
s_rom(282) <= -978;
s_rom(283) <= -974;
s_rom(284) <= -970;
s_rom(285) <= -965;
s_rom(286) <= -961;
s_rom(287) <= -956;
s_rom(288) <= -951;
s_rom(289) <= -945;
s_rom(290) <= -939;
s_rom(291) <= -933;
s_rom(292) <= -927;
s_rom(293) <= -920;
s_rom(294) <= -913;
s_rom(295) <= -906;
s_rom(296) <= -898;
s_rom(297) <= -891;
s_rom(298) <= -882;
s_rom(299) <= -874;
s_rom(300) <= -866;
s_rom(301) <= -857;
s_rom(302) <= -848;
s_rom(303) <= -838;
s_rom(304) <= -829;
s_rom(305) <= -819;
s_rom(306) <= -809;
s_rom(307) <= -798;
s_rom(308) <= -788;
s_rom(309) <= -777;
s_rom(310) <= -766;
s_rom(311) <= -754;
s_rom(312) <= -743;
s_rom(313) <= -731;
s_rom(314) <= -719;
s_rom(315) <= -707;
s_rom(316) <= -694;
s_rom(317) <= -681;
s_rom(318) <= -669;
s_rom(319) <= -656;
s_rom(320) <= -642;
s_rom(321) <= -629;
s_rom(322) <= -615;
s_rom(323) <= -601;
s_rom(324) <= -587;
s_rom(325) <= -573;
s_rom(326) <= -559;
s_rom(327) <= -544;
s_rom(328) <= -529;
s_rom(329) <= -515;
s_rom(330) <= -500;
s_rom(331) <= -484;
s_rom(332) <= -469;
s_rom(333) <= -453;
s_rom(334) <= -438;
s_rom(335) <= -422;
s_rom(336) <= -406;
s_rom(337) <= -390;
s_rom(338) <= -374;
s_rom(339) <= -358;
s_rom(340) <= -342;
s_rom(341) <= -325;
s_rom(342) <= -309;
s_rom(343) <= -292;
s_rom(344) <= -275;
s_rom(345) <= -258;
s_rom(346) <= -241;
s_rom(347) <= -224;
s_rom(348) <= -207;
s_rom(349) <= -190;
s_rom(350) <= -173;
s_rom(351) <= -156;
s_rom(352) <= -139;
s_rom(353) <= -121;
s_rom(354) <= -104;
s_rom(355) <= -87;
s_rom(356) <= -69;
s_rom(357) <= -52;
s_rom(358) <= -34;
s_rom(359) <= -17;
s_rom(360) <= 0;

c_rom(0) <= 1000;
c_rom(1) <= 999;
c_rom(2) <= 999;
c_rom(3) <= 998;
c_rom(4) <= 997;
c_rom(5) <= 996;
c_rom(6) <= 994;
c_rom(7) <= 992;
c_rom(8) <= 990;
c_rom(9) <= 987;
c_rom(10) <= 984;
c_rom(11) <= 981;
c_rom(12) <= 978;
c_rom(13) <= 974;
c_rom(14) <= 970;
c_rom(15) <= 965;
c_rom(16) <= 961;
c_rom(17) <= 956;
c_rom(18) <= 951;
c_rom(19) <= 945;
c_rom(20) <= 939;
c_rom(21) <= 933;
c_rom(22) <= 927;
c_rom(23) <= 920;
c_rom(24) <= 913;
c_rom(25) <= 906;
c_rom(26) <= 898;
c_rom(27) <= 891;
c_rom(28) <= 882;
c_rom(29) <= 874;
c_rom(30) <= 866;
c_rom(31) <= 857;
c_rom(32) <= 848;
c_rom(33) <= 838;
c_rom(34) <= 829;
c_rom(35) <= 819;
c_rom(36) <= 809;
c_rom(37) <= 798;
c_rom(38) <= 788;
c_rom(39) <= 777;
c_rom(40) <= 766;
c_rom(41) <= 754;
c_rom(42) <= 743;
c_rom(43) <= 731;
c_rom(44) <= 719;
c_rom(45) <= 707;
c_rom(46) <= 694;
c_rom(47) <= 681;
c_rom(48) <= 669;
c_rom(49) <= 656;
c_rom(50) <= 642;
c_rom(51) <= 629;
c_rom(52) <= 615;
c_rom(53) <= 601;
c_rom(54) <= 587;
c_rom(55) <= 573;
c_rom(56) <= 559;
c_rom(57) <= 544;
c_rom(58) <= 529;
c_rom(59) <= 515;
c_rom(60) <= 500;
c_rom(61) <= 484;
c_rom(62) <= 469;
c_rom(63) <= 453;
c_rom(64) <= 438;
c_rom(65) <= 422;
c_rom(66) <= 406;
c_rom(67) <= 390;
c_rom(68) <= 374;
c_rom(69) <= 358;
c_rom(70) <= 342;
c_rom(71) <= 325;
c_rom(72) <= 309;
c_rom(73) <= 292;
c_rom(74) <= 275;
c_rom(75) <= 258;
c_rom(76) <= 241;
c_rom(77) <= 224;
c_rom(78) <= 207;
c_rom(79) <= 190;
c_rom(80) <= 173;
c_rom(81) <= 156;
c_rom(82) <= 139;
c_rom(83) <= 121;
c_rom(84) <= 104;
c_rom(85) <= 87;
c_rom(86) <= 69;
c_rom(87) <= 52;
c_rom(88) <= 34;
c_rom(89) <= 17;
c_rom(90) <= 0;
c_rom(91) <= -17;
c_rom(92) <= -34;
c_rom(93) <= -52;
c_rom(94) <= -69;
c_rom(95) <= -87;
c_rom(96) <= -104;
c_rom(97) <= -121;
c_rom(98) <= -139;
c_rom(99) <= -156;
c_rom(100) <= -173;
c_rom(101) <= -190;
c_rom(102) <= -207;
c_rom(103) <= -224;
c_rom(104) <= -241;
c_rom(105) <= -258;
c_rom(106) <= -275;
c_rom(107) <= -292;
c_rom(108) <= -309;
c_rom(109) <= -325;
c_rom(110) <= -342;
c_rom(111) <= -358;
c_rom(112) <= -374;
c_rom(113) <= -390;
c_rom(114) <= -406;
c_rom(115) <= -422;
c_rom(116) <= -438;
c_rom(117) <= -453;
c_rom(118) <= -469;
c_rom(119) <= -484;
c_rom(120) <= -499;
c_rom(121) <= -515;
c_rom(122) <= -529;
c_rom(123) <= -544;
c_rom(124) <= -559;
c_rom(125) <= -573;
c_rom(126) <= -587;
c_rom(127) <= -601;
c_rom(128) <= -615;
c_rom(129) <= -629;
c_rom(130) <= -642;
c_rom(131) <= -656;
c_rom(132) <= -669;
c_rom(133) <= -681;
c_rom(134) <= -694;
c_rom(135) <= -707;
c_rom(136) <= -719;
c_rom(137) <= -731;
c_rom(138) <= -743;
c_rom(139) <= -754;
c_rom(140) <= -766;
c_rom(141) <= -777;
c_rom(142) <= -788;
c_rom(143) <= -798;
c_rom(144) <= -809;
c_rom(145) <= -819;
c_rom(146) <= -829;
c_rom(147) <= -838;
c_rom(148) <= -848;
c_rom(149) <= -857;
c_rom(150) <= -866;
c_rom(151) <= -874;
c_rom(152) <= -882;
c_rom(153) <= -891;
c_rom(154) <= -898;
c_rom(155) <= -906;
c_rom(156) <= -913;
c_rom(157) <= -920;
c_rom(158) <= -927;
c_rom(159) <= -933;
c_rom(160) <= -939;
c_rom(161) <= -945;
c_rom(162) <= -951;
c_rom(163) <= -956;
c_rom(164) <= -961;
c_rom(165) <= -965;
c_rom(166) <= -970;
c_rom(167) <= -974;
c_rom(168) <= -978;
c_rom(169) <= -981;
c_rom(170) <= -984;
c_rom(171) <= -987;
c_rom(172) <= -990;
c_rom(173) <= -992;
c_rom(174) <= -994;
c_rom(175) <= -996;
c_rom(176) <= -997;
c_rom(177) <= -998;
c_rom(178) <= -999;
c_rom(179) <= -999;
c_rom(180) <= -1000;
c_rom(181) <= -999;
c_rom(182) <= -999;
c_rom(183) <= -998;
c_rom(184) <= -997;
c_rom(185) <= -996;
c_rom(186) <= -994;
c_rom(187) <= -992;
c_rom(188) <= -990;
c_rom(189) <= -987;
c_rom(190) <= -984;
c_rom(191) <= -981;
c_rom(192) <= -978;
c_rom(193) <= -974;
c_rom(194) <= -970;
c_rom(195) <= -965;
c_rom(196) <= -961;
c_rom(197) <= -956;
c_rom(198) <= -951;
c_rom(199) <= -945;
c_rom(200) <= -939;
c_rom(201) <= -933;
c_rom(202) <= -927;
c_rom(203) <= -920;
c_rom(204) <= -913;
c_rom(205) <= -906;
c_rom(206) <= -898;
c_rom(207) <= -891;
c_rom(208) <= -882;
c_rom(209) <= -874;
c_rom(210) <= -866;
c_rom(211) <= -857;
c_rom(212) <= -848;
c_rom(213) <= -838;
c_rom(214) <= -829;
c_rom(215) <= -819;
c_rom(216) <= -809;
c_rom(217) <= -798;
c_rom(218) <= -788;
c_rom(219) <= -777;
c_rom(220) <= -766;
c_rom(221) <= -754;
c_rom(222) <= -743;
c_rom(223) <= -731;
c_rom(224) <= -719;
c_rom(225) <= -707;
c_rom(226) <= -694;
c_rom(227) <= -681;
c_rom(228) <= -669;
c_rom(229) <= -656;
c_rom(230) <= -642;
c_rom(231) <= -629;
c_rom(232) <= -615;
c_rom(233) <= -601;
c_rom(234) <= -587;
c_rom(235) <= -573;
c_rom(236) <= -559;
c_rom(237) <= -544;
c_rom(238) <= -529;
c_rom(239) <= -515;
c_rom(240) <= -500;
c_rom(241) <= -484;
c_rom(242) <= -469;
c_rom(243) <= -453;
c_rom(244) <= -438;
c_rom(245) <= -422;
c_rom(246) <= -406;
c_rom(247) <= -390;
c_rom(248) <= -374;
c_rom(249) <= -358;
c_rom(250) <= -342;
c_rom(251) <= -325;
c_rom(252) <= -309;
c_rom(253) <= -292;
c_rom(254) <= -275;
c_rom(255) <= -258;
c_rom(256) <= -241;
c_rom(257) <= -224;
c_rom(258) <= -207;
c_rom(259) <= -190;
c_rom(260) <= -173;
c_rom(261) <= -156;
c_rom(262) <= -139;
c_rom(263) <= -121;
c_rom(264) <= -104;
c_rom(265) <= -87;
c_rom(266) <= -69;
c_rom(267) <= -52;
c_rom(268) <= -34;
c_rom(269) <= -17;
c_rom(270) <= 0;
c_rom(271) <= 17;
c_rom(272) <= 34;
c_rom(273) <= 52;
c_rom(274) <= 69;
c_rom(275) <= 87;
c_rom(276) <= 104;
c_rom(277) <= 121;
c_rom(278) <= 139;
c_rom(279) <= 156;
c_rom(280) <= 173;
c_rom(281) <= 190;
c_rom(282) <= 207;
c_rom(283) <= 224;
c_rom(284) <= 241;
c_rom(285) <= 258;
c_rom(286) <= 275;
c_rom(287) <= 292;
c_rom(288) <= 309;
c_rom(289) <= 325;
c_rom(290) <= 342;
c_rom(291) <= 358;
c_rom(292) <= 374;
c_rom(293) <= 390;
c_rom(294) <= 406;
c_rom(295) <= 422;
c_rom(296) <= 438;
c_rom(297) <= 453;
c_rom(298) <= 469;
c_rom(299) <= 484;
c_rom(300) <= 500;
c_rom(301) <= 515;
c_rom(302) <= 529;
c_rom(303) <= 544;
c_rom(304) <= 559;
c_rom(305) <= 573;
c_rom(306) <= 587;
c_rom(307) <= 601;
c_rom(308) <= 615;
c_rom(309) <= 629;
c_rom(310) <= 642;
c_rom(311) <= 656;
c_rom(312) <= 669;
c_rom(313) <= 681;
c_rom(314) <= 694;
c_rom(315) <= 707;
c_rom(316) <= 719;
c_rom(317) <= 731;
c_rom(318) <= 743;
c_rom(319) <= 754;
c_rom(320) <= 766;
c_rom(321) <= 777;
c_rom(322) <= 788;
c_rom(323) <= 798;
c_rom(324) <= 809;
c_rom(325) <= 819;
c_rom(326) <= 829;
c_rom(327) <= 838;
c_rom(328) <= 848;
c_rom(329) <= 857;
c_rom(330) <= 866;
c_rom(331) <= 874;
c_rom(332) <= 882;
c_rom(333) <= 891;
c_rom(334) <= 898;
c_rom(335) <= 906;
c_rom(336) <= 913;
c_rom(337) <= 920;
c_rom(338) <= 927;
c_rom(339) <= 933;
c_rom(340) <= 939;
c_rom(341) <= 945;
c_rom(342) <= 951;
c_rom(343) <= 956;
c_rom(344) <= 961;
c_rom(345) <= 965;
c_rom(346) <= 970;
c_rom(347) <= 974;
c_rom(348) <= 978;
c_rom(349) <= 981;
c_rom(350) <= 984;
c_rom(351) <= 987;
c_rom(352) <= 990;
c_rom(353) <= 992;
c_rom(354) <= 994;
c_rom(355) <= 996;
c_rom(356) <= 997;
c_rom(357) <= 998;
c_rom(358) <= 999;
c_rom(359) <= 999;
c_rom(360) <= 1000;


            end if;
        end procedure rom_generator;
end package body fftpackage;